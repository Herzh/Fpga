module contador (ck, SQ);

	input ck;
	output [3:0